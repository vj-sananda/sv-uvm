package mypkg;
//import uvm_pkg::*;

`include "channel.svh"
typedef channel #(logic [8:0]) driver_channel ;

//`include "heartbeat.sv"

endpackage
  
