class ethernet_pkt extends uvm_transaction ;

rand byte preamble[8];

`uvm_object_utils(ethernet_pkt)

endclass
  
